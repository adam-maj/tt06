/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_adammaj (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
  alu alu_instance (
    .clk(clk),
    .reset(rst_n),
    .rs(ui_in[3:0]),
    .rt(ui_in[7:4]),
    .alu_arithmetic_mux(uio_in[1:0]),
    .alu_out(alu_out)
  );

  // All output pins must be assigned. If not used, assign to 0.
  assign uo_out  = {4'b0,alu_out};  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out = 0;
  assign uio_oe  = 0;
endmodule
